module ang_to_ascii (
    input wire [7:0] angle_in,
    output logic [11:0] ascii_out
);

always_comb begin
    case (angle_in)
        8'd0: ascii_out = 12'b000000000000;
        8'd1: ascii_out = 12'b000000000001;
        8'd2: ascii_out = 12'b000000000010;
        8'd3: ascii_out = 12'b000000000011;
        8'd4: ascii_out = 12'b000000000100;
        8'd5: ascii_out = 12'b000000000101;
        8'd6: ascii_out = 12'b000000000110;
        8'd7: ascii_out = 12'b000000000111;
        8'd8: ascii_out = 12'b000000001000;
        8'd9: ascii_out = 12'b000000001001;
        8'd10: ascii_out = 12'b000000010000;
        8'd11: ascii_out = 12'b000000010001;
        8'd12: ascii_out = 12'b000000010010;
        8'd13: ascii_out = 12'b000000010011;
        8'd14: ascii_out = 12'b000000010100;
        8'd15: ascii_out = 12'b000000010101;
        8'd16: ascii_out = 12'b000000010110;
        8'd17: ascii_out = 12'b000000010111;
        8'd18: ascii_out = 12'b000000011000;
        8'd19: ascii_out = 12'b000000011001;
        8'd20: ascii_out = 12'b000000100000;
        8'd21: ascii_out = 12'b000000100001;
        8'd22: ascii_out = 12'b000000100010;
        8'd23: ascii_out = 12'b000000100011;
        8'd24: ascii_out = 12'b000000100100;
        8'd25: ascii_out = 12'b000000100101;
        8'd26: ascii_out = 12'b000000100110;
        8'd27: ascii_out = 12'b000000100111;
        8'd28: ascii_out = 12'b000000101000;
        8'd29: ascii_out = 12'b000000101001;
        8'd30: ascii_out = 12'b000000110000;
        8'd31: ascii_out = 12'b000000110001;
        8'd32: ascii_out = 12'b000000110010;
        8'd33: ascii_out = 12'b000000110011;
        8'd34: ascii_out = 12'b000000110100;
        8'd35: ascii_out = 12'b000000110101;
        8'd36: ascii_out = 12'b000000110110;
        8'd37: ascii_out = 12'b000000110111;
        8'd38: ascii_out = 12'b000000111000;
        8'd39: ascii_out = 12'b000000111001;
        8'd40: ascii_out = 12'b000001000000;
        8'd41: ascii_out = 12'b000001000001;
        8'd42: ascii_out = 12'b000001000010;
        8'd43: ascii_out = 12'b000001000011;
        8'd44: ascii_out = 12'b000001000100;
        8'd45: ascii_out = 12'b000001000101;
        8'd46: ascii_out = 12'b000001000110;
        8'd47: ascii_out = 12'b000001000111;
        8'd48: ascii_out = 12'b000001001000;
        8'd49: ascii_out = 12'b000001001001;
        8'd50: ascii_out = 12'b000001010000;
        8'd51: ascii_out = 12'b000001010001;
        8'd52: ascii_out = 12'b000001010010;
        8'd53: ascii_out = 12'b000001010011;
        8'd54: ascii_out = 12'b000001010100;
        8'd55: ascii_out = 12'b000001010101;
        8'd56: ascii_out = 12'b000001010110;
        8'd57: ascii_out = 12'b000001010111;
        8'd58: ascii_out = 12'b000001011000;
        8'd59: ascii_out = 12'b000001011001;
        8'd60: ascii_out = 12'b000001100000;
        8'd61: ascii_out = 12'b000001100001;
        8'd62: ascii_out = 12'b000001100010;
        8'd63: ascii_out = 12'b000001100011;
        8'd64: ascii_out = 12'b000001100100;
        8'd65: ascii_out = 12'b000001100101;
        8'd66: ascii_out = 12'b000001100110;
        8'd67: ascii_out = 12'b000001100111;
        8'd68: ascii_out = 12'b000001101000;
        8'd69: ascii_out = 12'b000001101001;
        8'd70: ascii_out = 12'b000001110000;
        8'd71: ascii_out = 12'b000001110001;
        8'd72: ascii_out = 12'b000001110010;
        8'd73: ascii_out = 12'b000001110011;
        8'd74: ascii_out = 12'b000001110100;
        8'd75: ascii_out = 12'b000001110101;
        8'd76: ascii_out = 12'b000001110110;
        8'd77: ascii_out = 12'b000001110111;
        8'd78: ascii_out = 12'b000001111000;
        8'd79: ascii_out = 12'b000001111001;
        8'd80: ascii_out = 12'b000010000000;
        8'd81: ascii_out = 12'b000010000001;
        8'd82: ascii_out = 12'b000010000010;
        8'd83: ascii_out = 12'b000010000011;
        8'd84: ascii_out = 12'b000010000100;
        8'd85: ascii_out = 12'b000010000101;
        8'd86: ascii_out = 12'b000010000110;
        8'd87: ascii_out = 12'b000010000111;
        8'd88: ascii_out = 12'b000010001000;
        8'd89: ascii_out = 12'b000010001001;
        8'd90: ascii_out = 12'b000010010000;
        8'd91: ascii_out = 12'b000010010001;
        8'd92: ascii_out = 12'b000010010010;
        8'd93: ascii_out = 12'b000010010011;
        8'd94: ascii_out = 12'b000010010100;
        8'd95: ascii_out = 12'b000010010101;
        8'd96: ascii_out = 12'b000010010110;
        8'd97: ascii_out = 12'b000010010111;
        8'd98: ascii_out = 12'b000010011000;
        8'd99: ascii_out = 12'b000010011001;
        8'd100: ascii_out = 12'b000100000000;
        8'd101: ascii_out = 12'b000100000001;
        8'd102: ascii_out = 12'b000100000010;
        8'd103: ascii_out = 12'b000100000011;
        8'd104: ascii_out = 12'b000100000100;
        8'd105: ascii_out = 12'b000100000101;
        8'd106: ascii_out = 12'b000100000110;
        8'd107: ascii_out = 12'b000100000111;
        8'd108: ascii_out = 12'b000100001000;
        8'd109: ascii_out = 12'b000100001001;
        8'd110: ascii_out = 12'b000100010000;
        8'd111: ascii_out = 12'b000100010001;
        8'd112: ascii_out = 12'b000100010010;
        8'd113: ascii_out = 12'b000100010011;
        8'd114: ascii_out = 12'b000100010100;
        8'd115: ascii_out = 12'b000100010101;
        8'd116: ascii_out = 12'b000100010110;
        8'd117: ascii_out = 12'b000100010111;
        8'd118: ascii_out = 12'b000100011000;
        8'd119: ascii_out = 12'b000100011001;
        8'd120: ascii_out = 12'b000100100000;
        8'd121: ascii_out = 12'b000100100001;
        8'd122: ascii_out = 12'b000100100010;
        8'd123: ascii_out = 12'b000100100011;
        8'd124: ascii_out = 12'b000100100100;
        8'd125: ascii_out = 12'b000100100101;
        8'd126: ascii_out = 12'b000100100110;
        8'd127: ascii_out = 12'b000100100111;
        8'd128: ascii_out = 12'b000100101000;
        8'd129: ascii_out = 12'b000100101001;
        8'd130: ascii_out = 12'b000100110000;
        8'd131: ascii_out = 12'b000100110001;
        8'd132: ascii_out = 12'b000100110010;
        8'd133: ascii_out = 12'b000100110011;
        8'd134: ascii_out = 12'b000100110100;
        8'd135: ascii_out = 12'b000100110101;
        8'd136: ascii_out = 12'b000100110110;
        8'd137: ascii_out = 12'b000100110111;
        8'd138: ascii_out = 12'b000100111000;
        8'd139: ascii_out = 12'b000100111001;
        8'd140: ascii_out = 12'b000101000000;
        8'd141: ascii_out = 12'b000101000001;
        8'd142: ascii_out = 12'b000101000010;
        8'd143: ascii_out = 12'b000101000011;
        8'd144: ascii_out = 12'b000101000100;
        8'd145: ascii_out = 12'b000101000101;
        8'd146: ascii_out = 12'b000101000110;
        8'd147: ascii_out = 12'b000101000111;
        8'd148: ascii_out = 12'b000101001000;
        8'd149: ascii_out = 12'b000101001001;
        8'd150: ascii_out = 12'b000101010000;
        8'd151: ascii_out = 12'b000101010001;
        8'd152: ascii_out = 12'b000101010010;
        8'd153: ascii_out = 12'b000101010011;
        8'd154: ascii_out = 12'b000101010100;
        8'd155: ascii_out = 12'b000101010101;
        8'd156: ascii_out = 12'b000101010110;
        8'd157: ascii_out = 12'b000101010111;
        8'd158: ascii_out = 12'b000101011000;
        8'd159: ascii_out = 12'b000101011001;
        8'd160: ascii_out = 12'b000101100000;
        8'd161: ascii_out = 12'b000101100001;
        8'd162: ascii_out = 12'b000101100010;
        8'd163: ascii_out = 12'b000101100011;
        8'd164: ascii_out = 12'b000101100100;
        8'd165: ascii_out = 12'b000101100101;
        8'd166: ascii_out = 12'b000101100110;
        8'd167: ascii_out = 12'b000101100111;
        8'd168: ascii_out = 12'b000101101000;
        8'd169: ascii_out = 12'b000101101001;
        8'd170: ascii_out = 12'b000101110000;
        8'd171: ascii_out = 12'b000101110001;
        8'd172: ascii_out = 12'b000101110010;
        8'd173: ascii_out = 12'b000101110011;
        8'd174: ascii_out = 12'b000101110100;
        8'd175: ascii_out = 12'b000101110101;
        8'd176: ascii_out = 12'b000101110110;
        8'd177: ascii_out = 12'b000101110111;
        8'd178: ascii_out = 12'b000101111000;
        8'd179: ascii_out = 12'b000101111001;
        8'd180: ascii_out = 12'b000110000000;
        default: ascii_out = 0;
    endcase
end

endmodule